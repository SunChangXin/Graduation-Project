module seg_scan(
    input              clk         ,  // 系统时钟
    input              rst         ,  // 复位信号，高电平有效
    input      [2:0]   mode        ,  // 显示模式控制
    output reg [7:0]   row_sel     ,  // 行选择信号
    output reg [7:0]   col_sel     ,  // 列选择信号
    input      [63:0]  DianZhen_Data  // 显示数据，64位，控制8x8的数码管
);

	// 扫描频率和时钟频率的参数定义
	parameter   scanFreq   = 1250                       ;    // 扫描频率
	parameter   clkFreq    = 10000000                   ;    // 时钟频率  这两个参数很重要

	// 根据扫描频率和时钟频率计算扫描计数值
	parameter   cntNum  = clkFreq / (scanFreq * 8) - 1;

	reg[31:0]   scan_timer                                  ; // 扫描定时器
	reg[3:0]    scan_sel                                    ; // 扫描选择信号


	// 扫描定时器和扫描选择信号的控制逻辑
	always @(posedge clk or posedge rst)
	begin
		if(rst)
		begin
			scan_timer <= 32'd0;
			scan_sel <= 4'd0;
		end
		else if(scan_timer == cntNum)//>=
		begin
			scan_timer <= 32'd0;
			if(scan_sel == 4'd7)
				scan_sel <= 4'd0;
			else
				scan_sel <= scan_sel + 4'd1;
		end
		else
			begin
				scan_timer <= scan_timer + 32'd1;
			end
	end


	// 根据扫描选择信号和显示数据控制行列信号
	reg[7:0]    row_sel_reg                                 ; // 行选择寄存器
	reg[7:0]    col_sel_reg                                 ; // 列选择寄存器
	
	always@(*)//对每一行进行扫描
	begin
		case(scan_sel)
			4'd0://对第一行进行扫描
			begin
				col_sel_reg 			<= DianZhen_Data[(scan_sel+1)*8-1-:8]; //DianZhen_Data[7 -: 8] <–等价于–> DianZhen_Data[7:0]				
				row_sel_reg[7:1] 		<= 	7'b1111111;						
				if(DianZhen_Data[(scan_sel+1)*8-1-:8]>0)
				row_sel_reg[scan_sel]	<= 0;
				else
				row_sel_reg[scan_sel]	<= 1;
			end
			4'd1://对第二行进行扫描
			begin		
				col_sel_reg 			<= 	DianZhen_Data[(scan_sel+1)*8-1-:8];	//DianZhen_Data[15 -: 8] <–等价于–> DianZhen_Data[15:8]
				row_sel_reg[7:2] 		<= 	6'b111111;	
				row_sel_reg[0] 			<= 	1'b1;		
				
				if(DianZhen_Data[(scan_sel+1)*8-1-:8]>0)
				row_sel_reg[scan_sel]	<= 0;
				else
				row_sel_reg[scan_sel]	<= 1;
			end			
			4'd2://对第三行进行扫描
			begin
				col_sel_reg 			<= 	DianZhen_Data[(scan_sel+1)*8-1-:8];	//DianZhen_Data[23 -: 8] <–等价于–>DianZhen_Data[23:16]				
				row_sel_reg[7:3] 		<= 	5'b11111;		
				row_sel_reg[1:0] 		<= 	2'b11;					
				if(DianZhen_Data[(scan_sel+1)*8-1-:8]>0)
				row_sel_reg[scan_sel]	<= 0;
				else
				row_sel_reg[scan_sel]	<= 1;
			end
			4'd3://对第四行进行扫描
			begin
				col_sel_reg 			<= DianZhen_Data[(scan_sel+1)*8-1-:8];	//DianZhen_Data[31 -: 8] <–等价于–> DianZhen_Data[31:24]				
				row_sel_reg[7:4] 		<= 	4'b1111;		
				row_sel_reg[2:0] 		<= 	3'b111;		
				if(DianZhen_Data[(scan_sel+1)*8-1-:8]>0)
				row_sel_reg[scan_sel]	<= 0;
				else
				row_sel_reg[scan_sel]	<= 1;
			end
			4'd4://对第五行进行扫描
			begin
				col_sel_reg 			<= DianZhen_Data[(scan_sel+1)*8-1-:8];	//DianZhen_Data[39 -: 8] <–等价于–> DianZhen_Data[39:32]		
				
				row_sel_reg[7:5] 		<= 	3'b111;		
				row_sel_reg[3:0] 		<= 	4'b1111;				
				if(DianZhen_Data[(scan_sel+1)*8-1-:8]>0)
				row_sel_reg[scan_sel]	<= 0;
				else
				row_sel_reg[scan_sel]	<= 1;
			end
			4'd5://对第六行进行扫描
			begin
				col_sel_reg 			<= DianZhen_Data[(scan_sel+1)*8-1-:8];	//DianZhen_Data[47 -: 8] <–等价于–> DianZhen_Data[47:40]	
				row_sel_reg[7:6] 		<= 	2'b11;		
				row_sel_reg[4:0] 		<= 	5'b11111;					
				if(DianZhen_Data[(scan_sel+1)*8-1-:8]>0)
				row_sel_reg[scan_sel]	<= 0;
				else
				row_sel_reg[scan_sel]	<= 1;
			end
			4'd6://对第七行进行扫描                                                     //DianZhen_Data[55 -: 8] <–等价于–> DianZhen_Data[55:48]	
			begin
				col_sel_reg 			<= DianZhen_Data[(scan_sel+1)*8-1-:8];
				row_sel_reg[7] 			<= 	1'b1;		
				row_sel_reg[5:0] 		<= 	6'b111111;		

				if(DianZhen_Data[(scan_sel+1)*8-1-:8]>0)
				row_sel_reg[scan_sel]	<= 0;
				else
				row_sel_reg[scan_sel]	<= 1;
			end			
			4'd7: //对第八行进行扫描                                                    //DianZhen_Data[63 -: 8] <–等价于–> DianZhen_Data[63:56]
			begin	
				col_sel_reg 			<= DianZhen_Data[(scan_sel+1)*8-1-:8];			
				row_sel_reg[6:0] 		<= 	7'b1111111;	
				if(DianZhen_Data[(scan_sel+1)*8-1-:8]>0)
				row_sel_reg[scan_sel]	<= 0;
				else
				row_sel_reg[scan_sel]	<= 1;
			end						
			default:
			begin
				row_sel_reg <= 8'h00;
				col_sel_reg <= 8'h00;
			end
		endcase
	end
	

	always@(*)
	begin
		case(mode)       
			3'd1://左
				begin
					row_sel=row_sel_reg;
					col_sel={ col_sel_reg[0],col_sel_reg[1],col_sel_reg[2],col_sel_reg[3],col_sel_reg[4],col_sel_reg[5],col_sel_reg[6],col_sel_reg[7]};			
				end			

			3'd2://右
				begin
					 row_sel=row_sel_reg;
					 col_sel=col_sel_reg;			
				end
				
			3'd3://上
				begin
					row_sel=~{ col_sel_reg[0],col_sel_reg[1],col_sel_reg[2],col_sel_reg[3],col_sel_reg[4],col_sel_reg[5],col_sel_reg[6],col_sel_reg[7]};
					col_sel=~row_sel_reg;
				end					 
			
			3'd4://下	
				begin
					row_sel=~col_sel_reg;
					col_sel=~{row_sel_reg[0],row_sel_reg[1],row_sel_reg[2],row_sel_reg[3],row_sel_reg[4],row_sel_reg[5],row_sel_reg[6],row_sel_reg[7]};
				end					 				 
			
			default:
				begin
					row_sel=8'hff;
					col_sel=8'hff;	
				end
		endcase
	end
endmodule 