`timescale 1us / 1ns
module Counter_II_tb();
	
reg   clk;
reg   BTN0;
reg   BTN7;

wire  [7:0]  seg_sel;//(片选/位选)
wire  [7:0]  seg_led;//(段选)
wire  [7:0]  cout;


parameter CLK_PERIOD = 10;  //信号的定义，产生一个时钟信号j
always # (CLK_PERIOD/2)  clk = ~ clk;	

initial begin
	clk = 0;
	BTN0=1	;
	BTN7=1	;
	#2
	BTN0 = 0 ;	
	BTN7 = 0 ;		        //BTN7 = 1 ，解除复位
   
	#5000   press_BTN0;    //按一下BTN0键 暂停
   
	#5000   press_BTN0;    //按一下BTN0键 开始计数
	#10000   BTN7 = 1 ; //按下复位 清零
	#861000   press_BTN0;     //再按一下BTN0键 暂停

	#5000   press_BTN0;    //再按一下BTN0键 开始计数


	#10000   BTN7 = 1 ; //按下复位 清零

	#5000 	
	$stop;
end


Counter_II  u3 (
    .clk                     ( clk       ),
    .rst                     ( BTN7      ),
    .stop                    ( BTN0      ),
    .digtal_sw               ( seg_sel   ),
    .seg_led                 ( seg_led   ),
	 .count_out               ( cout      )
);

task press_BTN0;
	begin
			# (1*CLK_PERIOD )  BTN0 = 1; //抖动行为
			# (1*CLK_PERIOD )  BTN0 = 0; //抖动行为
			# (2*CLK_PERIOD )  BTN0 = 1; //抖动行为
			# (1*CLK_PERIOD )  BTN0 = 0; //抖动行为
			# (2*CLK_PERIOD )  BTN0 = 1; //抖动行为
			# (1*CLK_PERIOD )  BTN0 = 0; //抖动行为
			# (2*CLK_PERIOD )  BTN0 = 1; //抖动行为		
			# (10*CLK_PERIOD)  BTN0 = 1; //长时间的有效按键
			# (1*CLK_PERIOD )  BTN0 = 0;
		   #100;
	end
endtask


endmodule