module D_YM38(Ai,E1,E2_low,E3_low,ledx);
  
  input [3:0] Ai;
  input  E1;               //高电平有效使能端
  input  E2_low;           //低电平有效使能端
  input  E3_low;           //低电平有效使能
  
  reg a,b,c,d,e,f,g;
  reg [15:0] Y_low;
  
  
  output [6:0] ledx;
  
  
initial begin
  a <= 1'b0;
  b <= 1'b0;
  c <= 1'b0;
  d <= 1'b0;
  e <= 1'b0;
  f <= 1'b0;
  g <= 1'b0;
end  
  
always @ (Ai) begin
  if(E1 && ~E2_low && ~E3_low)
    case(Ai)
	 4'b0000: Y_low =16'b1111_1111_1111_1110;
	 4'b0001: Y_low =16'b1111_1111_1111_1101;
	 4'b0010: Y_low =16'b1111_1111_1111_1011;
	 4'b0011: Y_low =16'b1111_1111_1111_0111;
	 4'b0100: Y_low =16'b1111_1111_1110_1111;
	 4'b0101: Y_low =16'b1111_1111_1101_1111;
	 4'b0110: Y_low =16'b1111_1111_1011_1111;
	 4'b0111: Y_low =16'b1111_1111_0111_1111;
	 4'b1000: Y_low =16'b1111_1110_1111_1111;
	 4'b1001: Y_low =16'b1111_1101_1111_1111;
	 4'b1010: Y_low =16'b1111_1011_1111_1111;
	 4'b1011: Y_low =16'b1111_0111_1111_1111;
	 4'b1100: Y_low =16'b1110_1111_1111_1111;
	 4'b1101: Y_low =16'b1101_1111_1111_1111;
	 4'b1110: Y_low =16'b1011_1111_1111_1111;
	 4'b1111: Y_low =16'b0111_1111_1111_1111;
	 default: Y_low =16'b1111_1111_1111_1111;
    endcase 
  else
    Y_low =16'b1111_1111_1111_1111;
  
  if(!(Y[0] && Y[2] && Y[3] && Y[5] && Y[6] && Y[7] && Y[8] && Y[9]))
    a <= 1'b1;
	 
  if(!(Y[0] && Y[1] && Y[2] && Y[3] && Y[4] && Y[7] && Y[8] && Y[9]))
    b <= 1'b1;
	 
  if(!(Y[0] && Y[1] && Y[3] && Y[4] && Y[5] && Y[6] && Y[7] && Y[8] && Y[9]))
    c <= 1'b1;
	 
  if(!(Y[0] && Y[2] && Y[3] && Y[5] && Y[6] && Y[8] && Y[9]))
    d <= 1'b1;
	 
  if(!(Y[0] && Y[2] && Y[6] && Y[8]))
    e <= 1'b1;
	 
  if(!(Y[0] && Y[4] && Y[5] && Y[6] && Y[8] && Y[9]))
    f <= 1'b1;
	 
  if(!(Y[2] && Y[3] && Y[4] &&Y[5] && Y[6] && Y[8] && Y[9]))
    g <= 1'b1;
	 

  ledx = {a,b,c,d,e,f,g};
  
  
end  
  
  
  
  



endmodule