module StarT(BTN0);
	input BTN0;
	
	
	
	always @ (posedge BTN0)
	begin
		
		
		
		
	end
	
endmodule