module my_YiMa_7D(Ai,E1,E2_low,E3_low,ledx);
  
  input [3:0] Ai;
  input  E1;               //高电平有效使能端
  input  E2_low;           //低电平有效使能端
  input  E3_low;           //低电平有效使能
  
  reg a,b,c,d,e,f,g;
  reg [15:0] Y;
  
  
  output reg [6:0] ledx;
  
   
  
always @ (Ai or E1 or E2_low or E2_low) begin
  if(E1 && ~E2_low && ~E3_low)
    case(Ai)
	 4'b0000: Y =16'b1111_1111_1111_1110;
	 4'b0001: Y =16'b1111_1111_1111_1101;
	 4'b0010: Y =16'b1111_1111_1111_1011;
	 4'b0011: Y =16'b1111_1111_1111_0111;
	 4'b0100: Y =16'b1111_1111_1110_1111;
	 4'b0101: Y =16'b1111_1111_1101_1111;
	 4'b0110: Y =16'b1111_1111_1011_1111;
	 4'b0111: Y =16'b1111_1111_0111_1111;
	 4'b1000: Y =16'b1111_1110_1111_1111;
	 4'b1001: Y =16'b1111_1101_1111_1111;
	 4'b1010: Y =16'b1111_1011_1111_1111;
	 4'b1011: Y =16'b1111_0111_1111_1111;
	 4'b1100: Y =16'b1110_1111_1111_1111;
	 4'b1101: Y =16'b1101_1111_1111_1111;
	 4'b1110: Y =16'b1011_1111_1111_1111;
	 4'b1111: Y =16'b0111_1111_1111_1111;
	 default: Y =16'b1111_1111_1111_1111;
    endcase 
  else
    Y =16'b1111_1111_1111_1111;
  
  if(!(Y[0] && Y[2] && Y[3] && Y[5] && Y[6] && Y[7] && Y[8] && Y[9]))
    a <= 1'b1;
  if(Y[0] && Y[2] && Y[3] && Y[5] && Y[6] && Y[7] && Y[8] && Y[9])
    a <= 1'b0;
	 
  if(!(Y[0] && Y[1] && Y[2] && Y[3] && Y[4] && Y[7] && Y[8] && Y[9]))
    b <= 1'b1;
  if(Y[0] && Y[1] && Y[2] && Y[3] && Y[4] && Y[7] && Y[8] && Y[9])
    b <= 1'b0;
	 
  if(!(Y[0] && Y[1] && Y[3] && Y[4] && Y[5] && Y[6] && Y[7] && Y[8] && Y[9]))
    c <= 1'b1;
  if(Y[0] && Y[1] && Y[3] && Y[4] && Y[5] && Y[6] && Y[7] && Y[8] && Y[9])
    c <= 1'b0;
  
  if(!(Y[0] && Y[2] && Y[3] && Y[5] && Y[6] && Y[8] && Y[9]))
    d <= 1'b1;
  if(Y[0] && Y[2] && Y[3] && Y[5] && Y[6] && Y[8] && Y[9])
    d <= 1'b0;
  
  if(!(Y[0] && Y[2] && Y[6] && Y[8]))
    e <= 1'b1;
  if(Y[0] && Y[2] && Y[6] && Y[8])
    e <= 1'b0;
  
  if(!(Y[0] && Y[4] && Y[5] && Y[6] && Y[8] && Y[9]))
    f <= 1'b1;
  if(Y[0] && Y[4] && Y[5] && Y[6] && Y[8] && Y[9])
    f <= 1'b0;
  
  if(!(Y[2] && Y[3] && Y[4] &&Y[5] && Y[6] && Y[8] && Y[9]))
    g <= 1'b1;
  if(Y[2] && Y[3] && Y[4] &&Y[5] && Y[6] && Y[8] && Y[9])
    g <= 1'b0;
  

  ledx = {g,f,e,d,c,b,a};
  
  
end  
  
  
  
  



endmodule