module adder_1(a, b, Cin, Cout, Sum);
    input a, b, Cin;
	 output Cout, Sum;
	 wire x, y, z;
	 
	 
	 
	 xor xor1(x,a,b),
	     xor2(Sum,x,Cin);
	 and and1(y,a,b),
	     and2(z,Cin,x);
    or  or1(Cout,y,z);	 

endmodule
